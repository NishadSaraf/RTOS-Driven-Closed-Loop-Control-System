`timescale 1ns / 1ps

// n4fpga.v - Top level module for the ECE 544 Project - 2
//
// Copyright Chetan Bornarkar, Portland State University, 2016
// 
// Created By:	Roy Kravitz
// Modified By: Chetan Bornarkar
// Modified By: Nishad Saraf and Chaitanya Deshpande
// Date:		20-February-2017
// Version:		4.1
//
// Description:
// ------------
// This module provides the top level for the project 2 hardware.
// The module assume that PmodOLED and PmodHB3 are plugged into the JB and JA(bottom row) 
// expansion ports respectively and that a PmodENC is plugged into the JD expansion 
// port (bottom row).  
//////////////////////////////////////////////////////////////////////
module n4fpga(
    input				clk,			// 100Mhz clock input
    input				btnC,			// center pushbutton
    input				btnU,			// UP (North) pusbhbutton
    input				btnL,			// LEFT (West) pushbutton
    input				btnD,			// DOWN (South) pushbutton  - used for system reset
    input				btnR,			// RIGHT (East) pushbutton
	input				btnCpuReset,	// CPU reset pushbutton
    input	[15:0]		sw,				// slide switches on Nexys 4
    output	[15:0] 		led,			// LEDs on Nexys 4   
    output              RGB1_Blue,      // RGB1 LED (LD16) 
    output              RGB1_Green,
    output              RGB1_Red,
    output              RGB2_Blue,      // RGB2 LED (LD17)
    output              RGB2_Green,
    output              RGB2_Red,
    output [7:0]        an,             // Seven Segment display
    output [6:0]        seg,
    output              dp,             // decimal point display on the seven segment 
    
    input				uart_rtl_rxd,	// USB UART Rx and Tx on Nexys 4
    output				uart_rtl_txd,	
    
	inout   [7:0]       JA,             // JA PmodOLED connector 
	                                    // both rows are used 
    inout	[7:0] 		JB,				// JB Pmod connector 
                                        // Unused. Can be used for debuggin purposes 
    output	[7:0] 		JC,				// JC Pmod connector - debug signals
										// Can be used for debug purposes
	input	[7:0]		JD				// JD Pmod connector - PmodENC signals
);

// internal variables
// Clock and Reset 
wire				sysclk;              
wire				sysreset_n, sysreset;

// Rotary encoder 
wire				rotary_a, rotary_b, rotary_press, rotary_sw;

// PmodHB3
wire 	            HB3_DIR_OUT, HB3_EN, HB3_SA;

// GPIO pins 
//wire	[7:0]	    gpio_in;				// embsys GPIO input port
//wire	[7:0]	    gpio_out;				// embsys GPIO output port
wire    [4:0]       gpio_0_in;
wire    [15:0]      gpio_1_in;
//wire    [31:0]      gpio_2_in;
//wire    [15:0]      gpio_3_in;
wire    [15:0]      gpio_4_out;

// RGB LED 
wire                w_RGB1_Red, w_RGB1_Blue, w_RGB1_Green;

// LED pins 
wire    [15:0]      led_int;                // Nexys4IO drives these outputs

// Drive the leds from the signal generated by the microblaze 
//assign led = led_int;                   // LEDs are driven by led

// make the connections
// system-wide signals
assign sysclk = clk;
assign sysreset_n = btnCpuReset;		// The CPU reset pushbutton is asserted low.  The other pushbuttons are asserted high
										// but the microblaze for Nexys 4 expects reset to be asserted low
assign sysreset = ~sysreset_n;			// Generate a reset signal that is asserted high for any logic blocks expecting it.


// GPIO
assign gpio_0_in = {btnC,btnU,btnD,btnR,btnL};
assign led = gpio_4_out;

// PmodHB3 connections
assign JA[4] = HB3_DIR_OUT;
assign JA[5] = HB3_EN;
assign HB3_SA = JA[6]; 

// JC Connector pins can be used for debug purposes 
assign JC = 8'h00; 

// PmodENC signals
// JD - bottom row only
// Pins are assigned such that turning the knob to the right
// causes the rotary count to increment.
assign rotary_a = JD[5];
assign rotary_b = JD[4];
assign rotary_press = JD[6];
assign rotary_sw = JD[7];

// instantiate the embedded system
embsys EMBSYS
       (
	    // GPIO pins 
        .gpio_0_GPIO_tri_i(gpio_0_in),
        .gpio_1_GPIO_tri_i(sw),
        .gpio_4_GPIO_tri_o(gpio_4_out),
        //PMOD HB3 connections
        .PmodHB3_SA(HB3_SA),
        .PmodHB3_EN(HB3_EN),
        .PmodHB3_DIR(HB3_DIR_OUT),
        // Pmod Rotary Encoder
	    .pmodENC_A(rotary_a),
        .pmodENC_B(rotary_b),
        .pmodENC_btn(rotary_press),
        .pmodENC_sw(rotary_sw),
        // RGB1/2 Led's 
        .RGB1_Blue(RGB1_Blue),
        .RGB1_Green(RGB1_Green),
        .RGB1_Red(RGB1_Red),
        .RGB2_Blue(RGB2_Blue),
        .RGB2_Green(RGB2_Green),
        .RGB2_Red(RGB2_Red),
        // Seven Segment Display anode control  
        .an(an),
        .dp(dp),
        .led(led_int),
        .seg(seg),
        // Push buttons and switches  
        .btnC(btnC),
        .btnD(btnD),
        .btnL(btnL),
        .btnR(btnR),
        .btnU(btnU),
        .sw(sw),
        // reset and clock 
        .sysreset_n(sysreset_n),
        .sysclk(sysclk),
        // UART pins 
        .uart_rtl_rxd(uart_rtl_rxd),
        .uart_rtl_txd(uart_rtl_txd)
        );

endmodule